module snake_body(update,start,VGA_clk,snakeHead,snakeBody,xCount,yCount,x,y,z,w,h,size, data);
	input update , start,VGA_clk,xCount,yCount,x,y,w,z,h,size,data;
	wire[4:0] size ;
	wire reset ;
	output  snakeHead,snakeBody;
	reg [9:0] snakeX[0:31];
	reg [8:0] snakeY[0:31];
	reg [9:0] snakeHeadX;
	reg [9:0] snakeHeadY;
	integer  count1, count2, count3;
	reg snakeHead;
	reg snakeBody;
	wire [9:0] xCount;
	wire [9:0] yCount;
	wire [4:0] direction;
	wire displayArea;
	wire VGA_hSync, VGA_vSync, blank_n;
	wire [7:0] keyboard_data;
	
	Controller cont(x,y,z,w,h, direction, reset, VGA_clk);
	//kbInput k1(VGA_clk, data, direction, reset);
	//VGA_Controller1 (VGA_clk, xCount, yCount, displayArea, VGA_hSync, VGA_vSync, blank_n, keyboard_data, direction);
	
	always@(posedge update)
	begin
	if(start)
	begin
		if(direction != 5'b00111)begin
		for(count1 = 31; count1 > 0; count1 = count1 - 1)
			begin
				if(count1 <= size - 1)
				begin
					snakeX[count1] = snakeX[count1 - 1];
					snakeY[count1] = snakeY[count1 - 1];
				end
			end
			end
		case(direction)
			5'b00001: snakeY[0] <= (snakeY[0] - 10);
			5'b00010: snakeX[0] <= (snakeX[0] - 10);
			5'b00011: snakeY[0] <= (snakeY[0] + 10);
			5'b00100: snakeX[0] <= (snakeX[0] + 10);
			5'b00111:begin snakeX[0] <= snakeX[0];
			snakeY[0] <= snakeY[0]; end 
			endcase	
		end
	else if(~start)
	begin
		for(count3 = 1; count3 < 32; count3 = count3+1)
			begin
			snakeX[count3] = 700;
			snakeY[count3] = 500;
			end
			snakeX[0] = 300;
			snakeY[0] = 300;
	end
	
	end
	
	
	
	
	
	always@(posedge VGA_clk)
	begin
	
		snakeBody =0 ;
		
		for(count2 = 1; count2 < size; count2 = count2 + 1)
		begin
				
			if(snakeBody ==0 )
			snakeBody = ((xCount > snakeX[count2] && xCount < snakeX[count2]+10) && (yCount > snakeY[count2] && yCount < snakeY[count2]+10));
		
		
		end
	end


	
	always@(posedge VGA_clk)
	begin	
		snakeHead = (xCount > snakeX[0] && xCount < (snakeX[0]+10)) && (yCount > snakeY[0] && yCount < (snakeY[0]+10));
	end
	

endmodule 
